package packages;
    import uvm_pkg::*;

    // `include "sequence.svh"
    // `include "driver.svh"
    // `include "monitor.svh"
    // `include "agent.svh"
    // `include "scoreboard.svh"
    // `include "environment.svh"
    `include "test.svh"
endpackage