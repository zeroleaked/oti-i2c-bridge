`ifndef DUT_PARAMS_DEFINES
`define DUT_PARAMS_DEFINES

parameter DEFAULT_PRESCALE = 1;
parameter FIXED_PRESCALE = 0;
parameter CMD_FIFO = 1;
parameter CMD_FIFO_DEPTH = 32;
parameter WRITE_FIFO = 1;
parameter WRITE_FIFO_DEPTH = 32;
parameter READ_FIFO = 1;
parameter READ_FIFO_DEPTH = 32;

`endif