
`ifndef TIMESCALE_SV
`define TIMESCALE_SV
`timescale 1ns/1ps
`endif